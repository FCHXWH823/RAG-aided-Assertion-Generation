bind busarbiter busarbitersuit inst_busarbitersuit(.*); 