bind SEVEN SEVEN_sva #(.freq(freq), .CBITS(CBITS)) u_SEVEN_sva (.*);

