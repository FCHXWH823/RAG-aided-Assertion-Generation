bind simple_pipeline_en simple_pipeline_en_sva #(
    .WIDTH(WIDTH),
    .LATENCY(LATENCY)
    )
u_simple_pipeline_en_sva (.*);

