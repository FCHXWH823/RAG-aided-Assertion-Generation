bind rounding_division rounding_division_sva 
#(.DIV_LOG2(DIV_LOG2),
.OUT_WIDTH(OUT_WIDTH),
.IN_WIDTH(IN_WIDTH)) 
u_rounding_division_sva (.*);