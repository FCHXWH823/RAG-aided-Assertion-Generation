bind or1200_operandmuxes or1200_operandmuxes_sva #() u_or1200_operandmuxes_sva (.*);

