bind bit4counter bit4counter_sva #() u_bit4counter_sva (.*);

