bind a25_wishbone a25_wishbone_sva #() u_a25_wishbone_sva (.*);

