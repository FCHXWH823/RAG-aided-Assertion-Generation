bind Gray_To_Binary Gray_To_Binary_sva #(.DATA_WIDTH(DATA_WIDTH)) 
u_Gray_To_Binary_sva (.*);