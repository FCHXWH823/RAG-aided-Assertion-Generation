bind Flip_Flop_Array Flip_Flop_Array_sva 
#(.DATA_W(DATA_W),
  .ADDR_W(ADDR_W),
  .DATA_N(DATA_N)) 
u_Flip_Flop_Array_sva (.*);