
////////////////////////////////////////////////////////////////////////////////////////////////
////                                                              							////
////                                                              							////
////  	This file is part of the project                 									////
////	"instruction_list_pipelined_processor_with_peripherals"								////
////                                                              							////
////  http://opencores.org/project,instruction_list_pipelined_processor_with_peripherals	////
////                                                              							////
////                                                              							////
//// 				 Author:                                                  				////
////      			- Mahesh Sukhdeo Palve													////
////																						////
////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////
////																						////
//// 											                 							////
////                                                              							////
//// 					This source file may be used and distributed without         		////
//// 					restriction provided that this copyright statement is not    		////
//// 					removed from the file and that any derivative work contains  		////
//// 					the original copyright notice and the associated disclaimer. 		////
////                                                              							////
//// 					This source file is free software; you can redistribute it   		////
//// 					and/or modify it under the terms of the GNU Lesser General   		////
//// 					Public License as published by the Free Software Foundation; 		////
////					either version 2.1 of the License, or (at your option) any   		////
//// 					later version.                                               		////
////                                                             							////
//// 					This source is distributed in the hope that it will be       		////
//// 					useful, but WITHOUT ANY WARRANTY; without even the implied   		////
//// 					warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR      		////
//// 					PURPOSE.  See the GNU Lesser General Public License for more 		////
//// 					details.                                                     		////
////                                                              							////
//// 					You should have received a copy of the GNU Lesser General    		////
//// 					Public License along with this source; if not, download it   		////
//// 					from http://www.opencores.org/lgpl.shtml                     		////
////                                                              							////
////////////////////////////////////////////////////////////////////////////////////////////////

// 8-bit Pipelined Processor defines

`define		immDataLen			8

// program counter & instruction register
`define		instAddrLen			10			// 10-bit address => 1024 inst in rom
`define		instLen				15			// 15-bit fixed-length instructions
`define		instOpCodeLen		5
`define		instFieldLen		10


// control unit
`define		cuStateLen			4		// max 16 states
`define		END					`instOpCodeLen'b0
`define		JMP					`instOpCodeLen'b1
`define		Ld						`instOpCodeLen'b10
`define		Ldi					`instOpCodeLen'b11
`define		ST						`instOpCodeLen'b100
`define		ADD					`instOpCodeLen'b101
`define		SUB					`instOpCodeLen'b110
`define		MUL					`instOpCodeLen'b111
`define		DIV					`instOpCodeLen'b1000
`define		AND					`instOpCodeLen'b1001
`define		OR						`instOpCodeLen'b1010
`define		XOR					`instOpCodeLen'b1011
`define		GrT					`instOpCodeLen'b1100
`define		GE						`instOpCodeLen'b1101
`define		EQ						`instOpCodeLen'b1110
`define		LE						`instOpCodeLen'b1111
`define		LT						`instOpCodeLen'b10000
`define		PRE					`instOpCodeLen'b10001
`define		ETY					`instOpCodeLen'b10010
`define		RST					`instOpCodeLen'b10011
`define		LdTC					`instOpCodeLen'b10100
`define		LdACC					`instOpCodeLen'b10101
`define		UARTrd				`instOpCodeLen'b10110
`define		UARTwr				`instOpCodeLen'b10111
`define		UARTstat				`instOpCodeLen'b11000
//`define		SPIxFER				`instOpCodeLen'b11001
//`define		SPIstat				`instOpCodeLen'b11010
//`define		SPIwBUF				`instOpCodeLen'b11011
//`define		SPIrBUF				`instOpCodeLen'b11100

// alu opcodes
`define		aluOpcodeLen		4
`define		AND_alu				`aluOpcodeLen'b0
`define		OR_alu				`aluOpcodeLen'b1
`define		XOR_alu				`aluOpcodeLen'b10
`define		GT_alu				`aluOpcodeLen'b11
`define		GE_alu				`aluOpcodeLen'b100
`define		EQ_alu				`aluOpcodeLen'b101
`define		LE_alu				`aluOpcodeLen'b110
`define		LT_alu				`aluOpcodeLen'b111
`define		ADD_alu				`aluOpcodeLen'b1000
`define		SUB_alu				`aluOpcodeLen'b1001
`define		MUL_alu				`aluOpcodeLen'b1010
`define		DIV_alu				`aluOpcodeLen'b1011
`define		LD_data				`aluOpcodeLen'b1100

// bit RAM
`define		bitRamAddrLen		7		// 7-bit address
`define		bitRamDepth			128	// 2^7 = 128 locations

// byte RAM
`define		byteRamLen			8		// 8-bit input
`define		byteRamAddrLen		7		// 7-bit address
`define		byteRamDepth		128	// 2^7 = 128 locations

// input register
`define		inputNumber			128	// 128 inputs
`define		inputAddrLen		7		// 7-bit address

// output register
`define		outputNumber		128	// 128 outputs
`define		outputAddrLen		7		// 7-bit address

// accumulator multiplexer
`define		accMuxSelLen			4		// 2^4 = 16 selections available for accumulator
`define		accMuxSelImmData		`accMuxSelLen'b0
`define		accMuxSelAluOut		`accMuxSelLen'b1
`define		accMuxSelTcLoad		`accMuxSelLen'b10
`define		accMuxSelTcAcc			`accMuxSelLen'b11
`define		accMuxSelUartData		`accMuxSelLen'b100
`define		accMuxSelUartStat		`accMuxSelLen'b101

// operand2 multiplexer
`define		op2MuxSelLen			4		// 2^4 = 16 selections available for op2
`define		op2MuxSelInput			`op2MuxSelLen'b0
`define		op2MuxSelOutput		`op2MuxSelLen'b1
`define		op2MuxSelBitRam		`op2MuxSelLen'b10
`define		op2MuxSelByteRam		`op2MuxSelLen'b11
`define		op2MuxSel4			`op2MuxSelLen'b100
`define		op2MuxSel5			`op2MuxSelLen'b101
`define		op2MuxSel6			`op2MuxSelLen'b110

//-----------------------------------------------------------------------------------------------------

// peripheral defines
`define		timerAndCounter_peripheral
`define		UART_peripheral


//-----------------------------------------------------------------------------------------------------

// Timer-Counter
`define		tcAccLen				8		// 8-bit accumulated value
`define		tcPresetLen			8		// 8-bit preset value
`define		tcAddrLen			4
`define		tcTypeLen			2		// max 4-types
`define		tcNumbers			8		// total 8 modules (4-timers, 4-counters)

`define		timerType1			`tcTypeLen'b0
`define		timerType2			`tcTypeLen'b1
`define		timerType3			`tcTypeLen'b10

`define		counterType1		`tcTypeLen'b1
`define		counterType2		`tcTypeLen'b10


//-----------------------------------------------------------------------------------------------------

// UART
`define		dataBits 			8
`define		sbTick 				16	// ticks for stop bits (16 for 1-stopBit)
`define		fifoWidth 			4
`define 		number_fifo_regs 	16
`define 		fifoCntrWidth 		5
`define 		fifoDepth 			16

module bitRam_sva(
input reset,
input clk,
input bitRamEn,
input bitRamRw,
input bitRamIn,
input [`bitRamAddrLen-1:0] bitRamAddr,
input bitRamOut,
input bitRam [`bitRamDepth-1:0]
);

property a22;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[3] == 1 & bitRamAddr[4] == 1 & bitRamAddr[2] == 0) |-> (bitRamOut == 1);
endproperty
assert_a22: assert property(a22);

property a10;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[5] == 1 & bitRamAddr[3] == 0 & bitRamAddr[1] == 0) |-> (bitRamOut == 0);
endproperty
assert_a10: assert property(a10);

property a14;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[1] == 1 & bitRamAddr[2] == 0 & bitRamAddr[0] == 0 & bitRamAddr[3] == 0) |-> (bitRamOut == 0);
endproperty
assert_a14: assert property(a14);

property a16;
@(posedge clk) (bitRamRw == 1) ##1 (bitRamAddr[1] == 1 & bitRamAddr[2] == 1 & bitRamAddr[0] == 1 & bitRamAddr[5] == 1 & bitRamAddr[3] == 0) |-> (bitRamOut == 1);
endproperty
assert_a16: assert property(a16);

property a13;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[2] == 1 & bitRamAddr[1] == 0 & bitRamAddr[0] == 1 & bitRamAddr[4] == 0 & bitRamAddr[3] == 0) |-> (bitRamOut == 0);
endproperty
assert_a13: assert property(a13);

property a20;
@(posedge clk) (bitRamAddr[4] == 0 & bitRamAddr[2] == 0 & bitRamAddr[3] == 0 & bitRamAddr[5] == 0) |-> (bitRamOut == 1);
endproperty
assert_a20: assert property(a20);

property a17;
@(posedge clk) (bitRamAddr[2] == 0 & bitRamAddr[1] == 0 & bitRamAddr[3] == 0 & bitRamAddr[5] == 0) |-> (bitRamOut == 1);
endproperty
assert_a17: assert property(a17);

property a19;
@(posedge clk) (bitRamAddr[3] == 1 & bitRamAddr[1] == 1 & bitRamAddr[2] == 1 & bitRamAddr[0] == 1 & bitRamAddr[4] == 1 & bitRamAddr[5] == 1) |-> (bitRamOut == 1);
endproperty
assert_a19: assert property(a19);

property a9;
@(posedge clk) (bitRamAddr[0] == 0 & bitRamAddr[4] == 1 & bitRamAddr[1] == 0 & bitRamAddr[3] == 1 & bitRamAddr[2] == 0) |-> (bitRamOut == 0);
endproperty
assert_a9: assert property(a9);

property a21;
@(posedge clk) (bitRamRw == 1) ##1 (bitRamAddr[3] == 1 & bitRamIn == 0 & bitRamAddr[1] == 1 & bitRamAddr[0] == 0 & bitRamAddr[2] == 1) |-> (bitRamOut == 1);
endproperty
assert_a21: assert property(a21);

property a23;
@(posedge clk) (bitRamRw == 1) ##1 (bitRamAddr[3] == 1 & bitRamIn == 0 & bitRamAddr[1] == 1 & bitRamAddr[0] == 0 & bitRamAddr[4] == 0) |-> (bitRamOut == 1);
endproperty
assert_a23: assert property(a23);

property a25;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[4] == 0 & bitRamAddr[0] == 0 & bitRamIn == 0 & bitRamAddr[1] == 0 & bitRamAddr[2] == 1) |-> (bitRamOut == 1);
endproperty
assert_a25: assert property(a25);

property a29;
@(posedge clk) (bitRamRw == 1) ##1 (bitRamAddr[3] == 1 & bitRamIn == 0 & bitRamAddr[1] == 1 & bitRamAddr[4] == 1 & bitRamAddr[5] == 1) |-> (bitRamOut == 1);
endproperty
assert_a29: assert property(a29);

property a32;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[3] == 1 & bitRamAddr[4] == 1 & bitRamAddr[1] == 1 & bitRamIn == 0 & bitRamAddr[5] == 0) |-> (bitRamOut == 1);
endproperty
assert_a32: assert property(a32);

property a11;
@(posedge clk) (bitRamRw == 1) ##1 (bitRamAddr[2] == 1 & bitRamAddr[1] == 0 & bitRamIn == 1 & bitRamAddr[4] == 1 & bitRamAddr[0] == 1) |-> (bitRamOut == 0);
endproperty
assert_a11: assert property(a11);

property a6;
@(posedge clk) (bitRamRw == 1) ##1 (bitRamAddr[0] == 0 & bitRamAddr[4] == 1 & bitRamAddr[2] == 0 & bitRamIn == 0 & bitRamAddr[3] == 0) |-> (bitRamOut == 0);
endproperty
assert_a6: assert property(a6);

property a8;
@(posedge clk) (bitRamRw == 1) ##1 (bitRamAddr[5] == 0 & bitRamIn == 0 & bitRamAddr[4] == 0 & bitRamAddr[3] == 1 & bitRamAddr[0] == 1) |-> (bitRamOut == 0);
endproperty
assert_a8: assert property(a8);

property a24;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[3] == 1 & bitRamAddr[4] == 1 & bitRamIn == 1 & bitRamAddr[0] == 1) |-> (bitRamOut == 1);
endproperty
assert_a24: assert property(a24);

property a27;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[3] == 1 & bitRamIn == 0 & bitRamAddr[5] == 1 & bitRamAddr[0] == 1) |-> (bitRamOut == 1);
endproperty
assert_a27: assert property(a27);

property a33;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[3] == 1 & bitRamAddr[5] == 1 & bitRamAddr[4] == 1 & bitRamIn == 1) |-> (bitRamOut == 1);
endproperty
assert_a33: assert property(a33);

property a15;
@(posedge clk) (bitRamRw == 1) ##1 (bitRamAddr[1] == 1 & bitRamAddr[2] == 1 & bitRamAddr[0] == 1 & bitRamIn == 0) |-> (bitRamOut == 1);
endproperty
assert_a15: assert property(a15);

property a12;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[1] == 1 & bitRamIn == 1 & bitRamAddr[3] == 1 & bitRamAddr[4] == 0) |-> (bitRamOut == 0);
endproperty
assert_a12: assert property(a12);

property a1;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[1] == 0 & bitRamAddr[2] == 1 & bitRamIn == 1 & bitRamAddr[0] == 0) |-> (bitRamOut == 0);
endproperty
assert_a1: assert property(a1);

property a0;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[1] == 0 & bitRamAddr[2] == 1 & bitRamIn == 1 & bitRamAddr[3] == 0) |-> (bitRamOut == 0);
endproperty
assert_a0: assert property(a0);

property a28;
@(posedge clk) (bitRamAddr[4] == 0 & bitRamAddr[0] == 0 & bitRamIn == 0 & bitRamAddr[5] == 1 & bitRamAddr[1] == 0 & bitRamAddr[2] == 1 & bitRamAddr[3] == 0) |-> (bitRamOut == 1);
endproperty
assert_a28: assert property(a28);

property a30;
@(posedge clk) (bitRamAddr[3] == 1 & bitRamIn == 0 & bitRamAddr[5] == 1 & bitRamAddr[0] == 1 & bitRamAddr[1] == 0 & bitRamAddr[4] == 0) |-> (bitRamOut == 1);
endproperty
assert_a30: assert property(a30);

property a3;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[5] == 1 & bitRamIn == 1 & bitRamAddr[1] == 0) |-> (bitRamOut == 0);
endproperty
assert_a3: assert property(a3);

property a5;
@(posedge clk) (bitRamRw == 0) ##1 (bitRamAddr[5] == 1 & bitRamIn == 1 & bitRamAddr[2] == 0) |-> (bitRamOut == 0);
endproperty
assert_a5: assert property(a5);

property a26;
@(posedge clk) (bitRamAddr[4] == 0 & bitRamAddr[0] == 0 & bitRamAddr[2] == 0 & bitRamAddr[3] == 0 & bitRamIn == 1) |-> (bitRamOut == 1);
endproperty
assert_a26: assert property(a26);

property a31;
@(posedge clk) (bitRamAddr[1] == 1 & bitRamAddr[2] == 1 & bitRamAddr[5] == 0 & bitRamAddr[4] == 0 & bitRamIn == 1) |-> (bitRamOut == 1);
endproperty
assert_a31: assert property(a31);

property a18;
@(posedge clk) (bitRamAddr[3] == 1 & bitRamAddr[1] == 1 & bitRamIn == 0 & bitRamAddr[4] == 1 & bitRamAddr[0] == 1) |-> (bitRamOut == 1);
endproperty
assert_a18: assert property(a18);

property a2;
@(posedge clk) (bitRamAddr[1] == 0 & bitRamAddr[2] == 1 & bitRamIn == 1 & bitRamAddr[3] == 0 & bitRamAddr[0] == 0) |-> (bitRamOut == 0);
endproperty
assert_a2: assert property(a2);

property a4;
@(posedge clk) (bitRamAddr[1] == 0 & bitRamAddr[2] == 1 & bitRamIn == 1 & bitRamAddr[3] == 0 & bitRamAddr[4] == 1) |-> (bitRamOut == 0);
endproperty
assert_a4: assert property(a4);

property a7;
@(posedge clk) (bitRamAddr[1] == 0 & bitRamAddr[2] == 1 & bitRamIn == 1 & bitRamAddr[0] == 0 & bitRamAddr[4] == 0) |-> (bitRamOut == 0);
endproperty
assert_a7: assert property(a7);

endmodule