bind apb
 apb_sva u_apb_sva(
.PCLK(PCLK),
.TX_EMPTY(TX_EMPTY),
.INTERNAL_I2C_REGISTER_CONFIG(INTERNAL_I2C_REGISTER_CONFIG),
.RD_ENA(RD_ENA),
.READ_DATA_ON_RX(READ_DATA_ON_RX),
.PSELx(PSELx),
.INT_RX(INT_RX),
.WR_ENA(WR_ENA),
.INTERNAL_I2C_REGISTER_TIMEOUT(INTERNAL_I2C_REGISTER_TIMEOUT),
.RX_EMPTY(RX_EMPTY),
.INT_TX(INT_TX),
.ERROR(ERROR),
.PREADY(PREADY),
.PENABLE(PENABLE),
.PSLVERR(PSLVERR),
.PRESETn(PRESETn),
.PRDATA(PRDATA),
.PADDR(PADDR),
.WRITE_DATA_ON_TX(WRITE_DATA_ON_TX),
.PWRITE(PWRITE),
.PWDATA(PWDATA)
);