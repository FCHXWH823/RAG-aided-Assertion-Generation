bind simple_pipeline simple_pipeline_sva #(
    .WIDTH(WIDTH),
    .LATENCY(LATENCY)
    )
u_simple_pipeline_sva (.*);

