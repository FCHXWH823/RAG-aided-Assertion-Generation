bind i2c i2c_sva #(.divider(divider),.CBITS(CBITS)) u_i2c_sva (.*);

