
module module_i2c_sva(PCLK,PRESETn,fifo_tx_f_full,fifo_tx_f_empty,fifo_tx_data_out,fifo_rx_data_in,fifo_rx_f_full,fifo_rx_f_empty,fifo_rx_wr_en,
fifo_tx_rd_en,RX_EMPTY,TX_EMPTY,ERROR,ENABLE_SCL,ENABLE_SDA,SDA,SCL,DATA_CONFIG_REG,TIMEOUT_TX,state_tx,count_receive_data,RESPONSE,SDA_OUT,count_timeout,count_send_data,next_state_rx,BR_CLK_O,next_state_tx, count_tx,count_rx,BR_CLK_O_RX,SDA_OUT_RX,state_rx);

input PCLK;
input PRESETn;

//INTERFACE WITH FIFO TRANSMISSION
input fifo_tx_f_full;
input fifo_tx_f_empty;
input [32-1:0] fifo_tx_data_out;

//INTERFACE WITH FIFO RECEIVER
input fifo_rx_f_full;
input fifo_rx_f_empty;
input fifo_rx_wr_en;
input [32-1:0] fifo_rx_data_in; 

//INTERFACE WITH REGISTER CONFIGURATION
input [14-1:0] DATA_CONFIG_REG;
input [14-1:0] TIMEOUT_TX;

//INTERFACE TO APB AND READ FOR FIFO   
input fifo_tx_rd_en;
input   TX_EMPTY;
input   RX_EMPTY;
input ERROR;
input ENABLE_SDA;
input ENABLE_SCL;


//I2C BI DIRETIONAL PORTS
input SDA;
input SCL;
//registers
input state_tx;
input state_rx;
input count_receive_data;
input SDA_OUT;
input RESPONSE;
input count_timeout;
input count_send_data;
input next_state_rx;
input BR_CLK_O;
input next_state_tx;
input SDA_OUT_RX;
input count_tx;
input count_rx;
input BR_CLK_O_RX;

property a1;
@(posedge PCLK) (fifo_rx_f_empty == 1) |-> (RX_EMPTY == 1);
endproperty
assert_a1: assert property(a1);

property a0;
@(posedge PCLK) (fifo_rx_f_empty == 0) |-> (RX_EMPTY == 0);
endproperty
assert_a0: assert property(a0);

property a3;
@(posedge PCLK) (fifo_rx_f_empty == 1) |-> (RX_EMPTY == 1);
endproperty
assert_a3: assert property(a3);

property a2;
@(posedge PCLK) (fifo_rx_f_empty == 0) |-> (RX_EMPTY == 0);
endproperty
assert_a2: assert property(a2);

property a5;
@(posedge PCLK) (DATA_CONFIG_REG[1] == 0) |-> (ERROR == 0);
endproperty
assert_a5: assert property(a5);

property a4;
@(posedge PCLK) (DATA_CONFIG_REG[0] == 0) |-> (ERROR == 0);
endproperty
assert_a4: assert property(a4);

property a6;
@(posedge PCLK) (DATA_CONFIG_REG[0] == 1 & DATA_CONFIG_REG[1] == 1) |-> (ERROR == 1);
endproperty
assert_a6: assert property(a6);

endmodule