bind PWM PWM_sva #(.CBITS(CBITS)) u_PWM_sva (.*);

