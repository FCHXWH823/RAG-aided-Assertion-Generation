bind create_folder.sh create_folder.sh_sva #() u_create_folder.sh_sva (.*);

