bind register register_sva #(.WIDTH(WIDTH)) u_register_sva (.*);
