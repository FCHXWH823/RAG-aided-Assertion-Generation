bind PSGBusArb
 PSGBusArb_sva u_PSGBusArb_sva(
.rst(rst),
.ce(ce),
.sel2(sel2),
.sel4(sel4),
.req4(req4),
.req3(req3),
.req7(req7),
.clk(clk),
.sel1(sel1),
.sel0(sel0),
.seln(seln),
.sel3(sel3),
.ack(ack),
.req5(req5),
.req0(req0),
.sel6(sel6),
.sel5(sel5),
.req6(req6),
.sel7(sel7),
.req2(req2),
.req1(req1)
);