bind Gray_Code_Counter Gray_Code_Counter_sva #(.DATA_WIDTH(DATA_WIDTH)) 
u_Gray_Code_Counter_sva (.*);