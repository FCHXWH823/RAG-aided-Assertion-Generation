bind fpu_sub
 fpu_sub_sva u_fpu_sub_sva(
.mana_gtet_manb(mana_gtet_manb),
.fpu_op(fpu_op),
.subtra_shift(subtra_shift),
.diffshift_gt_exponent(diffshift_gt_exponent),
.mantissa_b(mantissa_b),
.large_norm_small_denorm(large_norm_small_denorm),
.diff(diff),
.opb(opb),
.subtra_shift_nonzero(subtra_shift_nonzero),
.exponent_large(exponent_large),
.in_norm_out_denorm(in_norm_out_denorm),
.diffshift_et_55(diffshift_et_55),
.clk(clk),
.rst(rst),
.enable(enable),
.minuend(minuend),
.small_is_denorm(small_is_denorm),
.expa_et_expb(expa_et_expb),
.exponent_2(exponent_2),
.exponent_small(exponent_small),
.diff_2(diff_2),
.sign(sign),
.subtra_shift_3(subtra_shift_3),
.a_gtet_b(a_gtet_b),
.mantissa_small(mantissa_small),
.subtra_shift_2(subtra_shift_2),
.subtrahend(subtrahend),
.diff_shift_2(diff_shift_2),
.opa(opa),
.expa_gt_expb(expa_gt_expb),
.small_is_nonzero(small_is_nonzero),
.exponent_b(exponent_b),
.exponent_a(exponent_a),
.mantissa_large(mantissa_large),
.diff_shift(diff_shift),
.mantissa_a(mantissa_a),
.exponent(exponent),
.exponent_diff(exponent_diff),
.diff_1(diff_1),
.subtra_fraction_enable(subtra_fraction_enable),
.large_is_denorm(large_is_denorm)
);