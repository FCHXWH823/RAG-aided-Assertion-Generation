bind control_unit control_unit_sva u_control_unit_sva(
      .sbox_sel(sbox_sel),
          .rk_sel(rk_sel),
          .key_out_sel(key_out_sel),
          .col_sel(col_sel),
          .key_en(key_en),
          .col_en(col_en),
         .round(round),
         .bypass_rk(bypass_rk),
         .bypass_key_en(bypass_key_en),
         .key_sel(key_sel),
         .iv_cnt_en(iv_cnt_en),
         .iv_cnt_sel(iv_cnt_sel),
         .key_derivation_en(key_derivation_en),
         .end_comp(end_comp),
         .key_init(key_init),
         .key_gen(key_gen),
         .mode_ctr(mode_ctr),
         .mode_cbc(mode_cbc),
         .last_round(last_round),
   	.encrypt_decrypt(encrypt_decrypt),
          .operation_mode(operation_mode),
          .aes_mode(aes_mode),
         .start(start),
         .disable_core(disable_core),
         .clk(clk),
         .rst_n(rst_n),
 .state(state), 
.next_state(next_state),
 .rd_count(rd_count),
.rd_count_en(rd_count_en),
 .op_key_derivation(op_key_derivation),
 .first_round(first_round),
 .op_mode(op_mode),
 .enc_dec(enc_dec)

);