
module control_unit_sva(
        input  [2:0] sbox_sel,
        input  [1:0] rk_sel,
        input  [1:0] key_out_sel,
        input  [1:0] col_sel,
        input  [3:0] key_en,
        input  [3:0] col_en,
        input  [3:0] round,
        input  bypass_rk,
        input  bypass_key_en,
        input  key_sel,
        input  iv_cnt_en,
        input  iv_cnt_sel,
        input  key_derivation_en,
        input end_comp,
        input key_init,
        input key_gen,
        input mode_ctr,
        input mode_cbc,
        input last_round,
  	input encrypt_decrypt,
        input [1:0] operation_mode,
        input [1:0] aes_mode,
        input start,
        input disable_core,
        input clk,
        input rst_n,
	input first_round,
	input state,
	input op_mode,
	input rd_count_en,
	input next_state,
	input rd_count,
	input op_key_derivation,
	input enc_dec
);
property a3;
@(posedge clk) (aes_mode[0] == 1) |-> (mode_ctr == 0);
endproperty
assert_a3: assert property(a3);

property a2;
@(posedge clk) (aes_mode[0] == 0) |-> (mode_cbc == 0);
endproperty
assert_a2: assert property(a2);

property a1;
@(posedge clk) (start == 0) |-> (key_init == 0);
endproperty
assert_a1: assert property(a1);

property a0;
@(posedge clk) (start == 1) |-> (key_init == 1);
endproperty
assert_a0: assert property(a0);

endmodule