bind gray gray_sva #(.CBITS(CBITS)) u_gray_sva (.*);

