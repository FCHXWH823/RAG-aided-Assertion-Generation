module arb2_sva(
input gnt1, gnt2,
input state,
input clk, rst,
input req1,
input req2
);


property a3;
@(posedge clk) (state == 1 & req2 == 1) |-> (gnt1 == 0);
endproperty
assert_a3: assert property(a3);

property a1;
@(posedge clk) (req1 == 1 & state == 0) |-> (gnt1 == 1);
endproperty
assert_a1: assert property(a1);

property a2;
@(posedge clk) (req1 == 0) |-> (gnt1 == 0);
endproperty
assert_a2: assert property(a2);

property a0;
@(posedge clk) (req1 == 1 & req2 == 0) |-> (gnt1 == 1);
endproperty
assert_a0: assert property(a0);

property a5;
@(posedge clk) (req1 == 1 & state == 0) |-> (gnt2 == 0);
endproperty
assert_a5: assert property(a5);

property a7;
@(posedge clk) (req2 == 1 & state == 1) |-> (gnt2 == 1);
endproperty
assert_a7: assert property(a7);

property a4;
@(posedge clk) (req2 == 0) |-> (gnt2 == 0);
endproperty
assert_a4: assert property(a4);

property a6;
@(posedge clk) (req2 == 1 & req1 == 0) |-> (gnt2 == 1);
endproperty
assert_a6: assert property(a6);

endmodule
