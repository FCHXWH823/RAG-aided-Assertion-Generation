bind counter counter_sva #(.MAX_AMOUNT(MAX_AMOUNT)) u_counter_sva (.*);

