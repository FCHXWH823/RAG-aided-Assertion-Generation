bind uart_transmit uart_transmit_sva #() u_uart_transmit_sva (.*);

