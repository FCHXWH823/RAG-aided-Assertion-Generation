bind lcd lcd_sva #(.clk_freq(clk_freq), .CBITS(CBITS)) u_lcd_sva (.*);

