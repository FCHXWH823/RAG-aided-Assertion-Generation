bind thermocouple thermocouple_sva u_thermocouple_sva (.*);

