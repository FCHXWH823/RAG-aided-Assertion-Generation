bind Ripple_Carry_Adder Ripple_Carry_Adder_sva #() u_Ripple_Carry_Adder_sva (.*);

