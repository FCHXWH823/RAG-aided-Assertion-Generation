bind simple_req_ack simple_req_ack_sva u_simple_req_ack_sva (.*);

