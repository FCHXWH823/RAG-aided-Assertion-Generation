bind Delay Delay_sva #(.N(N),.CBITS(CBITS)) u_Delay_sva (.*);

