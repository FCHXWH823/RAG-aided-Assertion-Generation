bind Programmable_Sequence_Detector Programmable_Sequence_Detector_sva #(.SEQ_W(SEQ_W)) 
u_Programmable_Sequence_Detector_sva (.*);