bind three_processor_bin_2 three_processor_bin_2_sva #() u_three_processor_bin_2_sva (.*);

