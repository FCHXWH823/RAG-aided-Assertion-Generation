bind AR AR_sva u_AR_sva (.*);

