bind simple_router simple_router_sva #(.DATA_WIDTH(DATA_WIDTH)) 
u_simple_router_sva(.*);