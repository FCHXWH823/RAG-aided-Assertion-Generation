module fifo_mem_sva#(parameter DEPTH=8, DATA_WIDTH=8, PTR_WIDTH=3)(
  input full, empty,
  input [PTR_WIDTH:0] b_wptr, b_rptr,
  input [DATA_WIDTH-1:0] fifo[0:DEPTH-1],
  input [DATA_WIDTH-1:0] data_out,
  input [DATA_WIDTH-1:0] data_in,
  input DEFAULT_CLOCK,
  input DEFAULT_RESET,
  input wclk, w_en, rclk, r_en
);

assert property(@(posedge DEFAULT_CLOCK) (w_en && !full) |-> (fifo[b_wptr[PTR_WIDTH-1:0]] == data_in));
assert property(@(posedge DEFAULT_CLOCK) (r_en && !empty) |-> (data_out == fifo[b_rptr[PTR_WIDTH-1:0]]));
assert property(@(posedge DEFAULT_CLOCK) (full) |-> (w_en == 0));
assert property(@(posedge DEFAULT_CLOCK) (empty) |-> (r_en == 0));
assert property(@(posedge DEFAULT_CLOCK) (w_en && full) |-> (fifo[b_wptr[PTR_WIDTH-1:0]] != data_in));
assert property(@(posedge DEFAULT_CLOCK) (r_en && empty) |-> (data_out == fifo[b_rptr[PTR_WIDTH-1:0]]));
assert property(@(posedge DEFAULT_CLOCK) (w_en && !full && r_en && !empty) |-> (fifo[b_wptr[PTR_WIDTH-1:0]] == data_in && data_out == fifo[b_rptr[PTR_WIDTH-1:0]]));
endmodule