bind Parallel_In_Serial_Out_Shift_Reg Parallel_In_Serial_Out_Shift_Reg_sva #(.DATA_WIDTH(DATA_WIDTH)) 
u_Parallel_In_Serial_Out_Shift_Reg_sva (.*);