bind host_interface
 host_interface_sva u_host_interface_sva(
.crc_init_en(crc_init_en),
.sample_bus(sample_bus),
.hwrite_pp(hwrite_pp),
.bus_wr(bus_wr),
.HWDATA(HWDATA),
.read_en(read_en),
.buffer_write_en(buffer_write_en),
.crc_init_out(crc_init_out),
.HSElx(HSElx),
.hsize_pp(hsize_pp),
.crc_cr_sel(crc_cr_sel),
.haddr_pp(haddr_pp),
.hselx_pp(hselx_pp),
.rev_out_type(rev_out_type),
.crc_cr_rd(crc_cr_rd),
.buffer_full(buffer_full),
.crc_idr_en(crc_idr_en),
.HCLK(HCLK),
.crc_cr_en(crc_cr_en),
.crc_poly_out(crc_poly_out),
.HADDR(HADDR),
.HSIZE(HSIZE),
.HREADYOUT(HREADYOUT),
.crc_init_sel(crc_init_sel),
.reset_chain(reset_chain),
.crc_idr_out(crc_idr_out),
.HTRANS(HTRANS),
.crc_poly_sel(crc_poly_sel),
.htrans_pp(htrans_pp),
.write_en(write_en),
.crc_poly_en(crc_poly_en),
.buffer_read_en(buffer_read_en),
.crc_out(crc_out),
.HRDATA(HRDATA),
.HWRITE(HWRITE),
.HREADY(HREADY),
.read_wait(read_wait),
.HRESETn(HRESETn),
.reset_pending(reset_pending),
.crc_dr_sel(crc_dr_sel),
.HRESP(HRESP),
.ahb_enable(ahb_enable),
.crc_cr_ff(crc_cr_ff),
.rev_in_type(rev_in_type),
.crc_poly_size(crc_poly_size),
.bus_size(bus_size),
.crc_idr_sel(crc_idr_sel)
);