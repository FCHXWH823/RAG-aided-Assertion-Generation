bind or1200_ctrl or1200_ctrl_sva #() u_or1200_ctrl_sva (.*);

