bind arbiter arbiter_sva #() u_arbiter_sva (.*);

