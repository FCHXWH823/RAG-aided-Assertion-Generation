bind reversing_bits reversing_bits_sva #(.DATA_WIDTH(DATA_WIDTH)) 
u_reversing_bits_sva (.*);