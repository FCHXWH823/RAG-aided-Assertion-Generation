bind ff ff_sva u_ff_sva (.*);
