bind or1200_if or1200_if_sva #() u_or1200_if_sva (.*);

