bind VGA VGA_sva #() u_VGA_sva (.*);

