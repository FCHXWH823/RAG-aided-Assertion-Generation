bind delay delay_sva #() u_delay_sva (.*);

