bind second_largest second_largest_sva #(.DATA_WIDTH(DATA_WIDTH)) 
u_second_largest_sva (.*);