bind module_i2c
 module_i2c_sva u_module_i2c_sva(
.PCLK(PCLK),
.RX_EMPTY(RX_EMPTY),
.fifo_tx_data_out(fifo_tx_data_out),
.count_rx(count_rx),
.BR_CLK_O_RX(BR_CLK_O_RX),
.ENABLE_SCL(ENABLE_SCL),
.SDA_OUT(SDA_OUT),
.PRESETn(PRESETn),
.state_rx(state_rx),
.fifo_rx_wr_en(fifo_rx_wr_en),
.RESPONSE(RESPONSE),
.BR_CLK_O(BR_CLK_O),
.count_receive_data(count_receive_data),
.SDA(SDA),
.count_send_data(count_send_data),
.DATA_CONFIG_REG(DATA_CONFIG_REG),
.TX_EMPTY(TX_EMPTY),
.count_timeout(count_timeout),
.TIMEOUT_TX(TIMEOUT_TX),
.ERROR(ERROR),
.SDA_OUT_RX(SDA_OUT_RX),
.fifo_rx_f_empty(fifo_rx_f_empty),
.state_tx(state_tx),
.SCL(SCL),
.fifo_rx_f_full(fifo_rx_f_full),
.fifo_tx_f_empty(fifo_tx_f_empty),
.count_tx(count_tx),
.ENABLE_SDA(ENABLE_SDA),
.fifo_rx_data_in(fifo_rx_data_in),
.next_state_rx(next_state_rx),
.next_state_tx(next_state_tx),
.fifo_tx_f_full(fifo_tx_f_full),
.fifo_tx_rd_en(fifo_tx_rd_en)
);